----------------------------------------------------------------------------------
-- CMS Muon Endcap
-- GEM Collaboration
-- Optohybrid v3 Firmware -- TDC
-- 2018/07/11 -- Initial
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

library work;
use work.types_pkg.all;
use work.param_pkg.all;
use work.ipbus_pkg.all;
use work.registers.all;

entity oh_tdc is
port(

    -- Clocks
    clk_1x_i : in std_logic;
    clk_8x_i : in std_logic;

    -- Config
    reset_i       : in std_logic;

    -- Inputs
    trigger_i   : in std_logic;
    sbits_i     : in std_logic_vector(23 downto 0);

    -- ipbus

    ipb_mosi_i : in  ipb_wbus;
    ipb_miso_o : out ipb_rbus;

    ipb_reset_i : in std_logic;
    ipb_clk_i : in std_logic

);
end oh_tdc;


architecture Behavioral of oh_tdc is

    signal reset : std_logic;
    signal reset_local : std_logic;
    signal resetting_o : std_logic;
    signal calibrate : std_logic;
    signal calibrating : std_logic;
    signal window_mask : std_logic_vector (255 downto 0);
    signal vfat_mask : std_logic_vector (23 downto 0);
    signal fifo_rden : std_logic_vector (23 downto 0);
    signal fifo_dout : std32_array_t (23 downto 0);
    signal fifo_valid : std_logic_vector (23 downto 0);
    signal fifo_underflow : std_logic_vector (23 downto 0);
    signal callut_addr : std_logic_vector(8 downto 0);
    signal callut_data : std_logic_vector(11 downto 0);

    ------ Register signals begin (this section is generated by <optohybrid_top>/tools/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_TDC_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_TDC_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_TDC_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_TDC_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_TDC_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_TDC_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_TDC_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_TDC_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_TDC_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------

begin

    process (clk_1x_i) begin
        if (rising_edge(clk_1x_i)) then
            reset <= reset_local or reset_i;
        end if;
    end process;

    tdc_inst : entity work.tdc
    port map (
        clk_1x_i => clk_1x_i,
        clk_8x_i => clk_8x_i,

        -- Config
        reset_i       => reset,
        resetting_o   => resetting_o,

        calibrate_i   => calibrate,
        calibrating_o => calibrating,

        window_mask_i => window_mask,
        vfat_mask_i   => vfat_mask,

        -- Inputs
        trigger_i  => trigger_i,
        sbits_i    => sbits_i,

        -- FIFOs
        fifo_rden      => fifo_rden,
        fifo_dout      => fifo_dout,
        fifo_valid     => fifo_valid,
        fifo_underflow => fifo_underflow,

        -- Calibration LUT
        callut_addr_i => callut_addr,
        callut_data_o => callut_data

    );

    --===============================================================================================
    -- (this section is generated by <optohybrid_top>/tools/generate_registers.py -- do not edit)
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_TDC_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_TDC_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_TDC_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => clk_1x_i,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"0";
    regs_addresses(1)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"1";
    regs_addresses(2)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"2";
    regs_addresses(3)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"3";
    regs_addresses(4)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"4";
    regs_addresses(5)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"5";
    regs_addresses(6)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"6";
    regs_addresses(7)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"7";
    regs_addresses(8)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"8";
    regs_addresses(9)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"9";
    regs_addresses(10)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"a";
    regs_addresses(11)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"b";
    regs_addresses(12)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"c";
    regs_addresses(13)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"d";
    regs_addresses(14)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"e";
    regs_addresses(15)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "00" & x"f";
    regs_addresses(16)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"0";
    regs_addresses(17)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"1";
    regs_addresses(18)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"2";
    regs_addresses(19)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"3";
    regs_addresses(20)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"4";
    regs_addresses(21)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"5";
    regs_addresses(22)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"6";
    regs_addresses(23)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"7";
    regs_addresses(24)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"8";
    regs_addresses(25)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"9";
    regs_addresses(26)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"a";
    regs_addresses(27)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"b";
    regs_addresses(28)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"c";
    regs_addresses(29)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"d";
    regs_addresses(30)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"e";
    regs_addresses(31)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "01" & x"f";
    regs_addresses(32)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"0";
    regs_addresses(33)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"1";
    regs_addresses(34)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"2";
    regs_addresses(35)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"3";
    regs_addresses(36)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"4";
    regs_addresses(37)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"5";
    regs_addresses(38)(REG_TDC_ADDRESS_MSB downto REG_TDC_ADDRESS_LSB) <= "10" & x"6";

    -- Connect read signals
    regs_read_arr(0)(REG_TDC_FIFO_rden_MSB downto REG_TDC_FIFO_rden_LSB) <= fifo_rden;
    regs_read_arr(1)(REG_TDC_FIFO_valid_MSB downto REG_TDC_FIFO_valid_LSB) <= fifo_valid;
    regs_read_arr(2)(REG_TDC_FIFO_underflow_MSB downto REG_TDC_FIFO_underflow_LSB) <= fifo_underflow;
    regs_read_arr(3)(REG_TDC_FIFO_dout0_MSB downto REG_TDC_FIFO_dout0_LSB) <= fifo_dout(0);
    regs_read_arr(4)(REG_TDC_FIFO_dout1_MSB downto REG_TDC_FIFO_dout1_LSB) <= fifo_dout(1);
    regs_read_arr(5)(REG_TDC_FIFO_dout2_MSB downto REG_TDC_FIFO_dout2_LSB) <= fifo_dout(2);
    regs_read_arr(6)(REG_TDC_FIFO_dout3_MSB downto REG_TDC_FIFO_dout3_LSB) <= fifo_dout(3);
    regs_read_arr(7)(REG_TDC_FIFO_dout4_MSB downto REG_TDC_FIFO_dout4_LSB) <= fifo_dout(4);
    regs_read_arr(8)(REG_TDC_FIFO_dout5_MSB downto REG_TDC_FIFO_dout5_LSB) <= fifo_dout(5);
    regs_read_arr(9)(REG_TDC_FIFO_dout6_MSB downto REG_TDC_FIFO_dout6_LSB) <= fifo_dout(6);
    regs_read_arr(10)(REG_TDC_FIFO_dout7_MSB downto REG_TDC_FIFO_dout7_LSB) <= fifo_dout(7);
    regs_read_arr(11)(REG_TDC_FIFO_dout8_MSB downto REG_TDC_FIFO_dout8_LSB) <= fifo_dout(8);
    regs_read_arr(12)(REG_TDC_FIFO_dout9_MSB downto REG_TDC_FIFO_dout9_LSB) <= fifo_dout(9);
    regs_read_arr(13)(REG_TDC_FIFO_dout10_MSB downto REG_TDC_FIFO_dout10_LSB) <= fifo_dout(10);
    regs_read_arr(14)(REG_TDC_FIFO_dout11_MSB downto REG_TDC_FIFO_dout11_LSB) <= fifo_dout(11);
    regs_read_arr(15)(REG_TDC_FIFO_dout12_MSB downto REG_TDC_FIFO_dout12_LSB) <= fifo_dout(12);
    regs_read_arr(16)(REG_TDC_FIFO_dout13_MSB downto REG_TDC_FIFO_dout13_LSB) <= fifo_dout(13);
    regs_read_arr(17)(REG_TDC_FIFO_dout14_MSB downto REG_TDC_FIFO_dout14_LSB) <= fifo_dout(14);
    regs_read_arr(18)(REG_TDC_FIFO_dout15_MSB downto REG_TDC_FIFO_dout15_LSB) <= fifo_dout(15);
    regs_read_arr(19)(REG_TDC_FIFO_dout16_MSB downto REG_TDC_FIFO_dout16_LSB) <= fifo_dout(16);
    regs_read_arr(20)(REG_TDC_FIFO_dout17_MSB downto REG_TDC_FIFO_dout17_LSB) <= fifo_dout(17);
    regs_read_arr(21)(REG_TDC_FIFO_dout18_MSB downto REG_TDC_FIFO_dout18_LSB) <= fifo_dout(18);
    regs_read_arr(22)(REG_TDC_FIFO_dout19_MSB downto REG_TDC_FIFO_dout19_LSB) <= fifo_dout(19);
    regs_read_arr(23)(REG_TDC_FIFO_dout20_MSB downto REG_TDC_FIFO_dout20_LSB) <= fifo_dout(20);
    regs_read_arr(24)(REG_TDC_FIFO_dout21_MSB downto REG_TDC_FIFO_dout21_LSB) <= fifo_dout(21);
    regs_read_arr(25)(REG_TDC_FIFO_dout22_MSB downto REG_TDC_FIFO_dout22_LSB) <= fifo_dout(22);
    regs_read_arr(26)(REG_TDC_FIFO_dout23_MSB downto REG_TDC_FIFO_dout23_LSB) <= fifo_dout(23);
    regs_read_arr(29)(REG_TDC_CTRL_CALIBRATING_BIT) <= calibrating;
    regs_read_arr(29)(REG_TDC_CTRL_CALLUT_DATA_MSB downto REG_TDC_CTRL_CALLUT_DATA_LSB) <= callut_data;
    regs_read_arr(29)(REG_TDC_CTRL_CALLUT_ADDR_MSB downto REG_TDC_CTRL_CALLUT_ADDR_LSB) <= callut_addr;
    regs_read_arr(30)(REG_TDC_CTRL_VFAT_MASK_MSB downto REG_TDC_CTRL_VFAT_MASK_LSB) <= vfat_mask;
    regs_read_arr(31)(REG_TDC_CTRL_WINDOW_MASK_0_MSB downto REG_TDC_CTRL_WINDOW_MASK_0_LSB) <= window_mask(31 downto 0);
    regs_read_arr(32)(REG_TDC_CTRL_WINDOW_MASK_1_MSB downto REG_TDC_CTRL_WINDOW_MASK_1_LSB) <= window_mask(63 downto 32);
    regs_read_arr(33)(REG_TDC_CTRL_WINDOW_MASK_2_MSB downto REG_TDC_CTRL_WINDOW_MASK_2_LSB) <= window_mask(95 downto 64);
    regs_read_arr(34)(REG_TDC_CTRL_WINDOW_MASK_3_MSB downto REG_TDC_CTRL_WINDOW_MASK_3_LSB) <= window_mask(127 downto 96);
    regs_read_arr(35)(REG_TDC_CTRL_WINDOW_MASK_4_MSB downto REG_TDC_CTRL_WINDOW_MASK_4_LSB) <= window_mask(159 downto 128);
    regs_read_arr(36)(REG_TDC_CTRL_WINDOW_MASK_5_MSB downto REG_TDC_CTRL_WINDOW_MASK_5_LSB) <= window_mask(191 downto 160);
    regs_read_arr(37)(REG_TDC_CTRL_WINDOW_MASK_6_MSB downto REG_TDC_CTRL_WINDOW_MASK_6_LSB) <= window_mask(223 downto 192);
    regs_read_arr(38)(REG_TDC_CTRL_WINDOW_MASK_7_MSB downto REG_TDC_CTRL_WINDOW_MASK_7_LSB) <= window_mask(255 downto 224);

    -- Connect write signals
    fifo_rden <= regs_write_arr(0)(REG_TDC_FIFO_rden_MSB downto REG_TDC_FIFO_rden_LSB);
    callut_addr <= regs_write_arr(29)(REG_TDC_CTRL_CALLUT_ADDR_MSB downto REG_TDC_CTRL_CALLUT_ADDR_LSB);
    vfat_mask <= regs_write_arr(30)(REG_TDC_CTRL_VFAT_MASK_MSB downto REG_TDC_CTRL_VFAT_MASK_LSB);
    window_mask(31 downto 0) <= regs_write_arr(31)(REG_TDC_CTRL_WINDOW_MASK_0_MSB downto REG_TDC_CTRL_WINDOW_MASK_0_LSB);
    window_mask(63 downto 32) <= regs_write_arr(32)(REG_TDC_CTRL_WINDOW_MASK_1_MSB downto REG_TDC_CTRL_WINDOW_MASK_1_LSB);
    window_mask(95 downto 64) <= regs_write_arr(33)(REG_TDC_CTRL_WINDOW_MASK_2_MSB downto REG_TDC_CTRL_WINDOW_MASK_2_LSB);
    window_mask(127 downto 96) <= regs_write_arr(34)(REG_TDC_CTRL_WINDOW_MASK_3_MSB downto REG_TDC_CTRL_WINDOW_MASK_3_LSB);
    window_mask(159 downto 128) <= regs_write_arr(35)(REG_TDC_CTRL_WINDOW_MASK_4_MSB downto REG_TDC_CTRL_WINDOW_MASK_4_LSB);
    window_mask(191 downto 160) <= regs_write_arr(36)(REG_TDC_CTRL_WINDOW_MASK_5_MSB downto REG_TDC_CTRL_WINDOW_MASK_5_LSB);
    window_mask(223 downto 192) <= regs_write_arr(37)(REG_TDC_CTRL_WINDOW_MASK_6_MSB downto REG_TDC_CTRL_WINDOW_MASK_6_LSB);
    window_mask(255 downto 224) <= regs_write_arr(38)(REG_TDC_CTRL_WINDOW_MASK_7_MSB downto REG_TDC_CTRL_WINDOW_MASK_7_LSB);

    -- Connect write pulse signals
    reset_local <= regs_write_pulse_arr(27);
    calibrate <= regs_write_pulse_arr(28);

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect counter instances

    -- Connect rate instances

    -- Connect read ready signals

    -- Defaults
    regs_defaults(0)(REG_TDC_FIFO_rden_MSB downto REG_TDC_FIFO_rden_LSB) <= REG_TDC_FIFO_rden_DEFAULT;
    regs_defaults(29)(REG_TDC_CTRL_CALLUT_ADDR_MSB downto REG_TDC_CTRL_CALLUT_ADDR_LSB) <= REG_TDC_CTRL_CALLUT_ADDR_DEFAULT;
    regs_defaults(30)(REG_TDC_CTRL_VFAT_MASK_MSB downto REG_TDC_CTRL_VFAT_MASK_LSB) <= REG_TDC_CTRL_VFAT_MASK_DEFAULT;
    regs_defaults(31)(REG_TDC_CTRL_WINDOW_MASK_0_MSB downto REG_TDC_CTRL_WINDOW_MASK_0_LSB) <= REG_TDC_CTRL_WINDOW_MASK_0_DEFAULT;
    regs_defaults(32)(REG_TDC_CTRL_WINDOW_MASK_1_MSB downto REG_TDC_CTRL_WINDOW_MASK_1_LSB) <= REG_TDC_CTRL_WINDOW_MASK_1_DEFAULT;
    regs_defaults(33)(REG_TDC_CTRL_WINDOW_MASK_2_MSB downto REG_TDC_CTRL_WINDOW_MASK_2_LSB) <= REG_TDC_CTRL_WINDOW_MASK_2_DEFAULT;
    regs_defaults(34)(REG_TDC_CTRL_WINDOW_MASK_3_MSB downto REG_TDC_CTRL_WINDOW_MASK_3_LSB) <= REG_TDC_CTRL_WINDOW_MASK_3_DEFAULT;
    regs_defaults(35)(REG_TDC_CTRL_WINDOW_MASK_4_MSB downto REG_TDC_CTRL_WINDOW_MASK_4_LSB) <= REG_TDC_CTRL_WINDOW_MASK_4_DEFAULT;
    regs_defaults(36)(REG_TDC_CTRL_WINDOW_MASK_5_MSB downto REG_TDC_CTRL_WINDOW_MASK_5_LSB) <= REG_TDC_CTRL_WINDOW_MASK_5_DEFAULT;
    regs_defaults(37)(REG_TDC_CTRL_WINDOW_MASK_6_MSB downto REG_TDC_CTRL_WINDOW_MASK_6_LSB) <= REG_TDC_CTRL_WINDOW_MASK_6_DEFAULT;
    regs_defaults(38)(REG_TDC_CTRL_WINDOW_MASK_7_MSB downto REG_TDC_CTRL_WINDOW_MASK_7_LSB) <= REG_TDC_CTRL_WINDOW_MASK_7_DEFAULT;

    -- Define writable regs
    regs_writable_arr(0) <= '1';
    regs_writable_arr(29) <= '1';
    regs_writable_arr(30) <= '1';
    regs_writable_arr(31) <= '1';
    regs_writable_arr(32) <= '1';
    regs_writable_arr(33) <= '1';
    regs_writable_arr(34) <= '1';
    regs_writable_arr(35) <= '1';
    regs_writable_arr(36) <= '1';
    regs_writable_arr(37) <= '1';
    regs_writable_arr(38) <= '1';

    --==== Registers end ============================================================================

end Behavioral;
