library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package sixbit_eightbit_pkg is

constant unused_key_0   : std_logic_vector (7 downto 0) := x"00"; -- 0b00000000 (disparity = -8)
constant unused_key_1   : std_logic_vector (7 downto 0) := x"01"; -- 0b00000001 (disparity = -6)
constant unused_key_2   : std_logic_vector (7 downto 0) := x"02"; -- 0b00000010 (disparity = -6)
constant unused_key_3   : std_logic_vector (7 downto 0) := x"03"; -- 0b00000011 (disparity = -4)
constant unused_key_4   : std_logic_vector (7 downto 0) := x"04"; -- 0b00000100 (disparity = -6)
constant unused_key_5   : std_logic_vector (7 downto 0) := x"05"; -- 0b00000101 (disparity = -4)
constant unused_key_6   : std_logic_vector (7 downto 0) := x"06"; -- 0b00000110 (disparity = -4)
constant unused_key_7   : std_logic_vector (7 downto 0) := x"07"; -- 0b00000111 (disparity = -2)
constant unused_key_8   : std_logic_vector (7 downto 0) := x"08"; -- 0b00001000 (disparity = -6)
constant unused_key_9   : std_logic_vector (7 downto 0) := x"09"; -- 0b00001001 (disparity = -4)
constant unused_key_10  : std_logic_vector (7 downto 0) := x"0A"; -- 0b00001010 (disparity = -4)
constant unused_key_11  : std_logic_vector (7 downto 0) := x"0B"; -- 0b00001011 (disparity = -2)
constant unused_key_12  : std_logic_vector (7 downto 0) := x"0C"; -- 0b00001100 (disparity = -4)
constant unused_key_13  : std_logic_vector (7 downto 0) := x"0D"; -- 0b00001101 (disparity = -2)
constant unused_key_14  : std_logic_vector (7 downto 0) := x"0E"; -- 0b00001110 (disparity = -2)
constant unused_key_15  : std_logic_vector (7 downto 0) := x"0F"; -- 0b00001111 (disparity = 0)
constant unused_key_16  : std_logic_vector (7 downto 0) := x"10"; -- 0b00010000 (disparity = -6)
constant unused_key_17  : std_logic_vector (7 downto 0) := x"11"; -- 0b00010001 (disparity = -4)
constant unused_key_18  : std_logic_vector (7 downto 0) := x"12"; -- 0b00010010 (disparity = -4)
constant unused_key_19  : std_logic_vector (7 downto 0) := x"13"; -- 0b00010011 (disparity = -2)
constant unused_key_20  : std_logic_vector (7 downto 0) := x"14"; -- 0b00010100 (disparity = -4)
constant unused_key_21  : std_logic_vector (7 downto 0) := x"15"; -- 0b00010101 (disparity = -2)
constant unused_key_22  : std_logic_vector (7 downto 0) := x"16"; -- 0b00010110 (disparity = -2)
constant unused_key_23  : std_logic_vector (7 downto 0) := x"18"; -- 0b00011000 (disparity = -4)
constant unused_key_24  : std_logic_vector (7 downto 0) := x"19"; -- 0b00011001 (disparity = -2)
constant unused_key_25  : std_logic_vector (7 downto 0) := x"1A"; -- 0b00011010 (disparity = -2)
constant unused_key_26  : std_logic_vector (7 downto 0) := x"1C"; -- 0b00011100 (disparity = -2)
constant unused_key_27  : std_logic_vector (7 downto 0) := x"1F"; -- 0b00011111 (disparity = 2)
constant unused_key_28  : std_logic_vector (7 downto 0) := x"20"; -- 0b00100000 (disparity = -6)
constant unused_key_29  : std_logic_vector (7 downto 0) := x"21"; -- 0b00100001 (disparity = -4)
constant unused_key_30  : std_logic_vector (7 downto 0) := x"22"; -- 0b00100010 (disparity = -4)
constant unused_key_31  : std_logic_vector (7 downto 0) := x"23"; -- 0b00100011 (disparity = -2)
constant unused_key_32  : std_logic_vector (7 downto 0) := x"24"; -- 0b00100100 (disparity = -4)
constant unused_key_33  : std_logic_vector (7 downto 0) := x"25"; -- 0b00100101 (disparity = -2)
constant unused_key_34  : std_logic_vector (7 downto 0) := x"26"; -- 0b00100110 (disparity = -2)
constant unused_key_35  : std_logic_vector (7 downto 0) := x"28"; -- 0b00101000 (disparity = -4)
constant unused_key_36  : std_logic_vector (7 downto 0) := x"29"; -- 0b00101001 (disparity = -2)
constant unused_key_37  : std_logic_vector (7 downto 0) := x"2A"; -- 0b00101010 (disparity = -2)
constant unused_key_38  : std_logic_vector (7 downto 0) := x"2C"; -- 0b00101100 (disparity = -2)
constant unused_key_39  : std_logic_vector (7 downto 0) := x"2F"; -- 0b00101111 (disparity = 2)
constant unused_key_40  : std_logic_vector (7 downto 0) := x"30"; -- 0b00110000 (disparity = -4)
constant unused_key_41  : std_logic_vector (7 downto 0) := x"31"; -- 0b00110001 (disparity = -2)
constant unused_key_42  : std_logic_vector (7 downto 0) := x"32"; -- 0b00110010 (disparity = -2)
constant unused_key_43  : std_logic_vector (7 downto 0) := x"34"; -- 0b00110100 (disparity = -2)
constant unused_key_44  : std_logic_vector (7 downto 0) := x"37"; -- 0b00110111 (disparity = 2)
constant unused_key_45  : std_logic_vector (7 downto 0) := x"38"; -- 0b00111000 (disparity = -2)
constant unused_key_46  : std_logic_vector (7 downto 0) := x"3B"; -- 0b00111011 (disparity = 2)
constant unused_key_47  : std_logic_vector (7 downto 0) := x"3D"; -- 0b00111101 (disparity = 2)
constant unused_key_48  : std_logic_vector (7 downto 0) := x"3E"; -- 0b00111110 (disparity = 2)
constant unused_key_49  : std_logic_vector (7 downto 0) := x"3F"; -- 0b00111111 (disparity = 4)
constant unused_key_50  : std_logic_vector (7 downto 0) := x"40"; -- 0b01000000 (disparity = -6)
constant unused_key_51  : std_logic_vector (7 downto 0) := x"41"; -- 0b01000001 (disparity = -4)
constant unused_key_52  : std_logic_vector (7 downto 0) := x"42"; -- 0b01000010 (disparity = -4)
constant unused_key_53  : std_logic_vector (7 downto 0) := x"43"; -- 0b01000011 (disparity = -2)
constant unused_key_54  : std_logic_vector (7 downto 0) := x"44"; -- 0b01000100 (disparity = -4)
constant unused_key_55  : std_logic_vector (7 downto 0) := x"45"; -- 0b01000101 (disparity = -2)
constant unused_key_56  : std_logic_vector (7 downto 0) := x"46"; -- 0b01000110 (disparity = -2)
constant unused_key_57  : std_logic_vector (7 downto 0) := x"47"; -- 0b01000111 (disparity = 0)
constant unused_key_58  : std_logic_vector (7 downto 0) := x"48"; -- 0b01001000 (disparity = -4)
constant unused_key_59  : std_logic_vector (7 downto 0) := x"49"; -- 0b01001001 (disparity = -2)
constant unused_key_60  : std_logic_vector (7 downto 0) := x"4A"; -- 0b01001010 (disparity = -2)
constant unused_key_61  : std_logic_vector (7 downto 0) := x"4C"; -- 0b01001100 (disparity = -2)
constant unused_key_62  : std_logic_vector (7 downto 0) := x"4F"; -- 0b01001111 (disparity = 2)
constant unused_key_63  : std_logic_vector (7 downto 0) := x"50"; -- 0b01010000 (disparity = -4)
constant unused_key_64  : std_logic_vector (7 downto 0) := x"51"; -- 0b01010001 (disparity = -2)
constant unused_key_65  : std_logic_vector (7 downto 0) := x"52"; -- 0b01010010 (disparity = -2)
constant unused_key_66  : std_logic_vector (7 downto 0) := x"54"; -- 0b01010100 (disparity = -2)
constant unused_key_67  : std_logic_vector (7 downto 0) := x"55"; -- 0b01010101 (disparity = 0)
constant unused_key_68  : std_logic_vector (7 downto 0) := x"57"; -- 0b01010111 (disparity = 2)
constant unused_key_69  : std_logic_vector (7 downto 0) := x"58"; -- 0b01011000 (disparity = -2)
constant unused_key_70  : std_logic_vector (7 downto 0) := x"5B"; -- 0b01011011 (disparity = 2)
constant unused_key_71  : std_logic_vector (7 downto 0) := x"5D"; -- 0b01011101 (disparity = 2)
constant unused_key_72  : std_logic_vector (7 downto 0) := x"5E"; -- 0b01011110 (disparity = 2)
constant unused_key_73  : std_logic_vector (7 downto 0) := x"5F"; -- 0b01011111 (disparity = 4)
constant unused_key_74  : std_logic_vector (7 downto 0) := x"60"; -- 0b01100000 (disparity = -4)
constant unused_key_75  : std_logic_vector (7 downto 0) := x"61"; -- 0b01100001 (disparity = -2)
constant unused_key_76  : std_logic_vector (7 downto 0) := x"62"; -- 0b01100010 (disparity = -2)
constant unused_key_77  : std_logic_vector (7 downto 0) := x"64"; -- 0b01100100 (disparity = -2)
constant unused_key_78  : std_logic_vector (7 downto 0) := x"67"; -- 0b01100111 (disparity = 2)
constant unused_key_79  : std_logic_vector (7 downto 0) := x"68"; -- 0b01101000 (disparity = -2)
constant unused_key_80  : std_logic_vector (7 downto 0) := x"6A"; -- 0b01101010 (disparity = 0)
constant unused_key_81  : std_logic_vector (7 downto 0) := x"6B"; -- 0b01101011 (disparity = 2)
constant unused_key_82  : std_logic_vector (7 downto 0) := x"6D"; -- 0b01101101 (disparity = 2)
constant unused_key_83  : std_logic_vector (7 downto 0) := x"6E"; -- 0b01101110 (disparity = 2)
constant unused_key_84  : std_logic_vector (7 downto 0) := x"6F"; -- 0b01101111 (disparity = 4)
constant unused_key_85  : std_logic_vector (7 downto 0) := x"70"; -- 0b01110000 (disparity = -2)
constant unused_key_86  : std_logic_vector (7 downto 0) := x"73"; -- 0b01110011 (disparity = 2)
constant unused_key_87  : std_logic_vector (7 downto 0) := x"75"; -- 0b01110101 (disparity = 2)
constant unused_key_88  : std_logic_vector (7 downto 0) := x"76"; -- 0b01110110 (disparity = 2)
constant unused_key_89  : std_logic_vector (7 downto 0) := x"77"; -- 0b01110111 (disparity = 4)
constant unused_key_90  : std_logic_vector (7 downto 0) := x"78"; -- 0b01111000 (disparity = 0)
constant unused_key_91  : std_logic_vector (7 downto 0) := x"79"; -- 0b01111001 (disparity = 2)
constant unused_key_92  : std_logic_vector (7 downto 0) := x"7A"; -- 0b01111010 (disparity = 2)
constant unused_key_93  : std_logic_vector (7 downto 0) := x"7B"; -- 0b01111011 (disparity = 4)
constant unused_key_94  : std_logic_vector (7 downto 0) := x"7C"; -- 0b01111100 (disparity = 2)
constant unused_key_95  : std_logic_vector (7 downto 0) := x"7D"; -- 0b01111101 (disparity = 4)
constant unused_key_96  : std_logic_vector (7 downto 0) := x"7E"; -- 0b01111110 (disparity = 4)
constant unused_key_97  : std_logic_vector (7 downto 0) := x"7F"; -- 0b01111111 (disparity = 6)
constant unused_key_98  : std_logic_vector (7 downto 0) := x"80"; -- 0b10000000 (disparity = -6)
constant unused_key_99  : std_logic_vector (7 downto 0) := x"81"; -- 0b10000001 (disparity = -4)
constant unused_key_100 : std_logic_vector (7 downto 0) := x"82"; -- 0b10000010 (disparity = -4)
constant unused_key_101 : std_logic_vector (7 downto 0) := x"83"; -- 0b10000011 (disparity = -2)
constant unused_key_102 : std_logic_vector (7 downto 0) := x"84"; -- 0b10000100 (disparity = -4)
constant unused_key_103 : std_logic_vector (7 downto 0) := x"85"; -- 0b10000101 (disparity = -2)
constant unused_key_104 : std_logic_vector (7 downto 0) := x"86"; -- 0b10000110 (disparity = -2)
constant unused_key_105 : std_logic_vector (7 downto 0) := x"88"; -- 0b10001000 (disparity = -4)
constant unused_key_106 : std_logic_vector (7 downto 0) := x"89"; -- 0b10001001 (disparity = -2)
constant unused_key_107 : std_logic_vector (7 downto 0) := x"8A"; -- 0b10001010 (disparity = -2)
constant unused_key_108 : std_logic_vector (7 downto 0) := x"8C"; -- 0b10001100 (disparity = -2)
constant unused_key_109 : std_logic_vector (7 downto 0) := x"8F"; -- 0b10001111 (disparity = 2)
constant unused_key_110 : std_logic_vector (7 downto 0) := x"90"; -- 0b10010000 (disparity = -4)
constant unused_key_111 : std_logic_vector (7 downto 0) := x"91"; -- 0b10010001 (disparity = -2)
constant unused_key_112 : std_logic_vector (7 downto 0) := x"92"; -- 0b10010010 (disparity = -2)
constant unused_key_113 : std_logic_vector (7 downto 0) := x"94"; -- 0b10010100 (disparity = -2)
constant unused_key_114 : std_logic_vector (7 downto 0) := x"97"; -- 0b10010111 (disparity = 2)
constant unused_key_115 : std_logic_vector (7 downto 0) := x"98"; -- 0b10011000 (disparity = -2)
constant unused_key_116 : std_logic_vector (7 downto 0) := x"9B"; -- 0b10011011 (disparity = 2)
constant unused_key_117 : std_logic_vector (7 downto 0) := x"9D"; -- 0b10011101 (disparity = 2)
constant unused_key_118 : std_logic_vector (7 downto 0) := x"9E"; -- 0b10011110 (disparity = 2)
constant unused_key_119 : std_logic_vector (7 downto 0) := x"9F"; -- 0b10011111 (disparity = 4)
constant unused_key_120 : std_logic_vector (7 downto 0) := x"A0"; -- 0b10100000 (disparity = -4)
constant unused_key_121 : std_logic_vector (7 downto 0) := x"A1"; -- 0b10100001 (disparity = -2)
constant unused_key_122 : std_logic_vector (7 downto 0) := x"A2"; -- 0b10100010 (disparity = -2)
constant unused_key_123 : std_logic_vector (7 downto 0) := x"A4"; -- 0b10100100 (disparity = -2)
constant unused_key_124 : std_logic_vector (7 downto 0) := x"A7"; -- 0b10100111 (disparity = 2)
constant unused_key_125 : std_logic_vector (7 downto 0) := x"A8"; -- 0b10101000 (disparity = -2)
constant unused_key_126 : std_logic_vector (7 downto 0) := x"AB"; -- 0b10101011 (disparity = 2)
constant unused_key_127 : std_logic_vector (7 downto 0) := x"AD"; -- 0b10101101 (disparity = 2)
constant unused_key_128 : std_logic_vector (7 downto 0) := x"AE"; -- 0b10101110 (disparity = 2)
constant unused_key_129 : std_logic_vector (7 downto 0) := x"AF"; -- 0b10101111 (disparity = 4)
constant unused_key_130 : std_logic_vector (7 downto 0) := x"B0"; -- 0b10110000 (disparity = -2)
constant unused_key_131 : std_logic_vector (7 downto 0) := x"B3"; -- 0b10110011 (disparity = 2)
constant unused_key_132 : std_logic_vector (7 downto 0) := x"B5"; -- 0b10110101 (disparity = 2)
constant unused_key_133 : std_logic_vector (7 downto 0) := x"B6"; -- 0b10110110 (disparity = 2)
constant unused_key_134 : std_logic_vector (7 downto 0) := x"B7"; -- 0b10110111 (disparity = 4)
constant unused_key_135 : std_logic_vector (7 downto 0) := x"B9"; -- 0b10111001 (disparity = 2)
constant unused_key_136 : std_logic_vector (7 downto 0) := x"BA"; -- 0b10111010 (disparity = 2)
constant unused_key_137 : std_logic_vector (7 downto 0) := x"BB"; -- 0b10111011 (disparity = 4)
constant unused_key_138 : std_logic_vector (7 downto 0) := x"BC"; -- 0b10111100 (disparity = 2)
constant unused_key_139 : std_logic_vector (7 downto 0) := x"BD"; -- 0b10111101 (disparity = 4)
constant unused_key_140 : std_logic_vector (7 downto 0) := x"BE"; -- 0b10111110 (disparity = 4)
constant unused_key_141 : std_logic_vector (7 downto 0) := x"BF"; -- 0b10111111 (disparity = 6)
constant unused_key_142 : std_logic_vector (7 downto 0) := x"C0"; -- 0b11000000 (disparity = -4)
constant unused_key_143 : std_logic_vector (7 downto 0) := x"C1"; -- 0b11000001 (disparity = -2)
constant unused_key_144 : std_logic_vector (7 downto 0) := x"C2"; -- 0b11000010 (disparity = -2)
constant unused_key_145 : std_logic_vector (7 downto 0) := x"C4"; -- 0b11000100 (disparity = -2)
constant unused_key_146 : std_logic_vector (7 downto 0) := x"C7"; -- 0b11000111 (disparity = 2)
constant unused_key_147 : std_logic_vector (7 downto 0) := x"C8"; -- 0b11001000 (disparity = -2)
constant unused_key_148 : std_logic_vector (7 downto 0) := x"CB"; -- 0b11001011 (disparity = 2)
constant unused_key_149 : std_logic_vector (7 downto 0) := x"CD"; -- 0b11001101 (disparity = 2)
constant unused_key_150 : std_logic_vector (7 downto 0) := x"CE"; -- 0b11001110 (disparity = 2)
constant unused_key_151 : std_logic_vector (7 downto 0) := x"CF"; -- 0b11001111 (disparity = 4)
constant unused_key_152 : std_logic_vector (7 downto 0) := x"D0"; -- 0b11010000 (disparity = -2)
constant unused_key_153 : std_logic_vector (7 downto 0) := x"D3"; -- 0b11010011 (disparity = 2)
constant unused_key_154 : std_logic_vector (7 downto 0) := x"D5"; -- 0b11010101 (disparity = 2)
constant unused_key_155 : std_logic_vector (7 downto 0) := x"D6"; -- 0b11010110 (disparity = 2)
constant unused_key_156 : std_logic_vector (7 downto 0) := x"D7"; -- 0b11010111 (disparity = 4)
constant unused_key_157 : std_logic_vector (7 downto 0) := x"D9"; -- 0b11011001 (disparity = 2)
constant unused_key_158 : std_logic_vector (7 downto 0) := x"DA"; -- 0b11011010 (disparity = 2)
constant unused_key_159 : std_logic_vector (7 downto 0) := x"DB"; -- 0b11011011 (disparity = 4)
constant unused_key_160 : std_logic_vector (7 downto 0) := x"DC"; -- 0b11011100 (disparity = 2)
constant unused_key_161 : std_logic_vector (7 downto 0) := x"DD"; -- 0b11011101 (disparity = 4)
constant unused_key_162 : std_logic_vector (7 downto 0) := x"DE"; -- 0b11011110 (disparity = 4)
constant unused_key_163 : std_logic_vector (7 downto 0) := x"DF"; -- 0b11011111 (disparity = 6)
constant unused_key_164 : std_logic_vector (7 downto 0) := x"E0"; -- 0b11100000 (disparity = -2)
constant unused_key_165 : std_logic_vector (7 downto 0) := x"E3"; -- 0b11100011 (disparity = 2)
constant unused_key_166 : std_logic_vector (7 downto 0) := x"E5"; -- 0b11100101 (disparity = 2)
constant unused_key_167 : std_logic_vector (7 downto 0) := x"E6"; -- 0b11100110 (disparity = 2)
constant unused_key_168 : std_logic_vector (7 downto 0) := x"E7"; -- 0b11100111 (disparity = 4)
constant unused_key_169 : std_logic_vector (7 downto 0) := x"E9"; -- 0b11101001 (disparity = 2)
constant unused_key_170 : std_logic_vector (7 downto 0) := x"EA"; -- 0b11101010 (disparity = 2)
constant unused_key_171 : std_logic_vector (7 downto 0) := x"EB"; -- 0b11101011 (disparity = 4)
constant unused_key_172 : std_logic_vector (7 downto 0) := x"EC"; -- 0b11101100 (disparity = 2)
constant unused_key_173 : std_logic_vector (7 downto 0) := x"ED"; -- 0b11101101 (disparity = 4)
constant unused_key_174 : std_logic_vector (7 downto 0) := x"EE"; -- 0b11101110 (disparity = 4)
constant unused_key_175 : std_logic_vector (7 downto 0) := x"EF"; -- 0b11101111 (disparity = 6)
constant unused_key_176 : std_logic_vector (7 downto 0) := x"F0"; -- 0b11110000 (disparity = 0)
constant unused_key_177 : std_logic_vector (7 downto 0) := x"F1"; -- 0b11110001 (disparity = 2)
constant unused_key_178 : std_logic_vector (7 downto 0) := x"F2"; -- 0b11110010 (disparity = 2)
constant unused_key_179 : std_logic_vector (7 downto 0) := x"F3"; -- 0b11110011 (disparity = 4)
constant unused_key_180 : std_logic_vector (7 downto 0) := x"F4"; -- 0b11110100 (disparity = 2)
constant unused_key_181 : std_logic_vector (7 downto 0) := x"F5"; -- 0b11110101 (disparity = 4)
constant unused_key_182 : std_logic_vector (7 downto 0) := x"F6"; -- 0b11110110 (disparity = 4)
constant unused_key_183 : std_logic_vector (7 downto 0) := x"F7"; -- 0b11110111 (disparity = 6)
constant unused_key_184 : std_logic_vector (7 downto 0) := x"F8"; -- 0b11111000 (disparity = 2)
constant unused_key_185 : std_logic_vector (7 downto 0) := x"F9"; -- 0b11111001 (disparity = 4)
constant unused_key_186 : std_logic_vector (7 downto 0) := x"FA"; -- 0b11111010 (disparity = 4)
constant unused_key_187 : std_logic_vector (7 downto 0) := x"FB"; -- 0b11111011 (disparity = 6)
constant unused_key_188 : std_logic_vector (7 downto 0) := x"FC"; -- 0b11111100 (disparity = 4)
constant unused_key_189 : std_logic_vector (7 downto 0) := x"FD"; -- 0b11111101 (disparity = 6)
constant unused_key_190 : std_logic_vector (7 downto 0) := x"FE"; -- 0b11111110 (disparity = 6)
constant unused_key_191 : std_logic_vector (7 downto 0) := x"FF"; -- 0b11111111 (disparity = 8)

constant IDLE_CHAR      : std_logic_vector (7 downto 0) := unused_key_69;
constant L1A_CHAR       : std_logic_vector (7 downto 0) := unused_key_80;
constant BC0_CHAR       : std_logic_vector (7 downto 0) := unused_key_159;
constant RESYNC_CHAR    : std_logic_vector (7 downto 0) := unused_key_136;

end sixbit_eightbit_pkg;
