----------------------------------------------------------------------------------
-- Company:        IIHE - ULB
-- Engineer:       Thomas Lenzi (thomas.lenzi@cern.ch)
-- 
-- Create Date:    11:22:49 06/30/2015 
-- Design Name:    OptoHybrid v2
-- Module Name:    vfat2_i2c_base - Behavioral 
-- Project Name:   OptoHybrid v2
-- Target Devices: xc6vlx130t-1ff1156
-- Tool versions:  ISE  P.20131013
-- Description: 
--
-- Handles I2C communications with the VFAT2
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity vfat2_i2c_base is
generic(
    CLK_DIV             : integer := 400
);
port(

    clk_i               : in std_logic;
    reset_i             : in std_logic;
    
    i2c_en_i            : in std_logic;
    i2c_address_i       : in std_logic_vector(6 downto 0);
    i2c_rw_i            : in std_logic;
    i2c_data_i          : in std_logic_vector(7 downto 0);
    
    i2c_valid_o         : out std_logic;
    i2c_error_o         : out std_logic;
    i2c_data_o          : out std_logic_vector(7 downto 0);
    
    vfat2_scl_o         : out std_logic;
    vfat2_sda_miso_i    : in std_logic;
    vfat2_sda_mosi_o    : out std_logic;
    vfat2_sda_tri_o     : out std_logic
    
);
end vfat2_i2c_base;

architecture Behavioral of vfat2_i2c_base is
    
    type state_t is (IDLE, START, ADDR, RW, RST_0, ACK_0, RD, ACK_1, RST_1, WR, RST_2, ACK_2, STOP, ERROR);
    
    signal state            : state_t;
    
    signal clk_divider      : integer range 0 to CLK_DIV;
    signal high_clk_pulse   : std_logic;
    signal low_clk_pulse    : std_logic;
    
    signal address          : std_logic_vector(6 downto 0);
    signal rw_n             : std_logic;
    signal din              : std_logic_vector(7 downto 0);
    signal dout             : std_logic_vector(7 downto 0);
    
    signal address_cnt      : integer range 0 to 6;
    signal data_cnt         : integer range 0 to 7;

begin

    --=========--
    --== SCK ==--
    --=========--
    
    process(clk_i)
    begin
        if (rising_edge(clk_i)) then
            if (reset_i = '1') then
                vfat2_scl_o <= '0';
                clk_divider <= 0;
                high_clk_pulse <= '0';
                low_clk_pulse <= '0';
            else
                -- Counting
                if (clk_divider = (CLK_DIV - 1)) then
                    clk_divider <= 0;
                else
                    clk_divider <= clk_divider + 1;
                end if;
                -- SCK generation
                if (clk_divider < (CLK_DIV - 1) / 2) then
                    vfat2_scl_o <= '1';
                else
                    vfat2_scl_o <= '0';
                end if;
                -- Start / Stop pulse & Read pulse
                if (clk_divider = (CLK_DIV - 1) / 4) then
                    high_clk_pulse <= '1';
                else
                    high_clk_pulse <= '0';
                end if;
                -- Data pulse
                if (clk_divider = (CLK_DIV - 1) * 3 / 4) then
                    low_clk_pulse <= '1';
                else
                    low_clk_pulse <= '0';
                end if;
            end if;
        end if;
    end process;

    --=========--
    --== SDA ==--
    --=========--

    process(clk_i)
    begin    
        if (rising_edge(clk_i)) then
            if (reset_i = '1') then
                vfat2_sda_mosi_o <= '1';
                vfat2_sda_tri_o <= '1';
                i2c_valid_o <= '0';
                i2c_error_o <= '0';
                i2c_data_o <= (others => '0');
                state <= IDLE;
            else
                case state is
                    -- IDLE
                    when IDLE =>
                        vfat2_sda_mosi_o <= '1';
                        vfat2_sda_tri_o <= '0';
                        i2c_valid_o <= '0';
                        i2c_error_o <= '0';
                        if (i2c_en_i = '1') then
                            state <= START;
                            address <= i2c_address_i;
                            rw_n <= i2c_rw_i;
                            din <= i2c_data_i;
                        end if;
                    -- Start
                    when START =>
                        if (high_clk_pulse = '1') then
                            vfat2_sda_mosi_o <= '0';
                            vfat2_sda_tri_o <= '0';
                            state <= ADDR;
                            address_cnt <= 6;
                        end if;
                    -- Address
                    when ADDR => 
                        if (low_clk_pulse = '1') then
                            vfat2_sda_mosi_o <= address(address_cnt);
                            vfat2_sda_tri_o <= '0';
                            if (address_cnt = 0) then
                                state <= RW;
                            else
                                address_cnt <= address_cnt - 1;
                            end if;
                        end if;
                    -- RW bit
                    when RW => 
                        if (low_clk_pulse = '1') then
                            vfat2_sda_mosi_o <= rw_n;
                            vfat2_sda_tri_o <= '0';
                            state <= RST_0;
                        end if;
                    -- Wait
                    when RST_0 => 
                        if (low_clk_pulse = '1') then
                            vfat2_sda_mosi_o <= '1';
                            vfat2_sda_tri_o <= '1';
                            state <= ACK_0;
                        end if;
                    -- Ackownledgment
                    when ACK_0 =>
                        if (high_clk_pulse = '1') then
                            vfat2_sda_mosi_o <= '1';
                            vfat2_sda_tri_o <= '1';
                            if (vfat2_sda_miso_i = '1') then
                                data_cnt <= 7;
                                case rw_n is
                                    when '1' => state <= RD;
                                    when others => state <= WR;
                                end case;
                            else
                                state <= ERROR;
                            end if;
                        end if;
                    -- Read
                    when RD => 
                        if (high_clk_pulse = '1') then
                            dout(data_cnt) <= vfat2_sda_miso_i;
                            vfat2_sda_mosi_o <= '1';
                            vfat2_sda_tri_o <= '1';
                            if (data_cnt = 7) then
                                state <= ACK_1;
                            else
                                data_cnt <= data_cnt - 1;
                            end if;
                        end if;
                    -- Read Ackownledgment 
                    when ACK_1 => 
                        if (low_clk_pulse = '1') then
                            vfat2_sda_mosi_o <= '1';
                            vfat2_sda_tri_o <= '0';
                            state <= RST_1;
                        end if;
                    -- Wait
                    when RST_1 => 
                        if (high_clk_pulse = '1') then
                            vfat2_sda_mosi_o <= '1';
                            vfat2_sda_tri_o <= '0';
                            state <= STOP;
                        end if;
                    -- Write
                    when WR => 
                        if (low_clk_pulse = '1') then
                            vfat2_sda_mosi_o <= dout(data_cnt);
                            vfat2_sda_tri_o <= '0';
                            if (data_cnt = 7) then
                                state <= RST_2;
                            else
                                data_cnt <= data_cnt - 1;
                            end if;
                        end if;
                    -- Wait
                    when RST_2 => 
                        if (low_clk_pulse = '1') then
                            vfat2_sda_mosi_o <= '1';
                            vfat2_sda_tri_o <= '1';
                            state <= ACK_2;
                        end if;
                    -- Write Ackownledgment 
                    when ACK_2 => 
                        if (high_clk_pulse = '1') then
                            vfat2_sda_mosi_o <= '1';
                            vfat2_sda_tri_o <= '1';
                            if (vfat2_sda_miso_i = '1') then
                                state <= STOP;
                            else
                                state <= ERROR;
                            end if;
                        end if;
                    -- STOP
                    when STOP => 
                        if (high_clk_pulse = '1') then
                            vfat2_sda_mosi_o <= '1';
                            vfat2_sda_tri_o <= '0';
                            i2c_valid_o <= '1';
                            i2c_error_o <= '0';
                            case rw_n is
                                when '1' => i2c_data_o <= dout;
                                when others => i2c_data_o <= (others => '0');
                            end case;
                            state <= IDLE;
                        end if;
                    -- ERROR
                    when ERROR => 
                        if (high_clk_pulse = '1') then
                            vfat2_sda_mosi_o <= '1';
                            vfat2_sda_tri_o <= '0';
                            i2c_valid_o <= '0';
                            i2c_error_o <= '1';
                            i2c_data_o <= (others => '0');
                            state <= IDLE;
                        end if;
                    --
                    when others => 
                        vfat2_sda_mosi_o <= '1';
                        vfat2_sda_tri_o <= '1';
                        i2c_valid_o <= '0';
                        i2c_error_o <= '0';
                        i2c_data_o <= (others => '0');
                        state <= IDLE;
                end case;  
            end if;
        end if;
    end process;
    
end Behavioral;