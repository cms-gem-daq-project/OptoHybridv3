
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package generation_pkg is
    constant RELEASE_HARDWARE       : std_logic_vector(7 downto  0) := x"2A";
end generation_pkg;
