----------------------------------------------------------------------------------
-- CMS Muon Endcap
-- GEM Collaboration
-- Optohybrid v3 Firmware -- Tap Delays
-- A. Peck
----------------------------------------------------------------------------------
-- Description:
--   This module holds trig polarity swaps derived from the Optohybrid PCB
----------------------------------------------------------------------------------
-- 2017/11/06 -- Initial
-- 2017/11/13 -- Port to vhdl
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package trig_pkg is

  constant DDR : integer := 0;
  constant MXSBITS : integer := 64 * (DDR+1);
  constant MXSBITS_CHAMBER : integer := 24*MXSBITS;

  constant  SOT_INVERT  : std_logic_vector (23 downto 0) :=
    '0' & -- SOF_INVERT[23]
    '1' & -- SOF_INVERT[22]
    '1' & -- SOF_INVERT[21]
    '0' & -- SOF_INVERT[20]
    '0' & -- SOF_INVERT[19]
    '1' & -- SOF_INVERT[18]
    '0' & -- SOF_INVERT[17]
    '1' & -- SOF_INVERT[16]
    '0' & -- SOF_INVERT[15]
    '1' & -- SOF_INVERT[14]
    '0' & -- SOF_INVERT[13]
    '0' & -- SOF_INVERT[12]
    '1' & -- SOF_INVERT[11]
    '0' & -- SOF_INVERT[10]
    '0' & -- SOF_INVERT[9]
    '1' & -- SOF_INVERT[8]
    '1' & -- SOF_INVERT[7]
    '0' & -- SOF_INVERT[6]
    '0' & -- SOF_INVERT[5]
    '1' & -- SOF_INVERT[4]
    '1' & -- SOF_INVERT[3]
    '1' & -- SOF_INVERT[2]
    '1' & -- SOF_INVERT[1]
    '1' ; -- SOF_INVERT[0]



  constant  TU_INVERT  : std_logic_vector (191 downto 0) :=
    '1' & -- TU_INVERT[191]
    '1' & -- TU_INVERT[190]
    '1' & -- TU_INVERT[189]
    '1' & -- TU_INVERT[188]
    '1' & -- TU_INVERT[187]
    '1' & -- TU_INVERT[186]
    '1' & -- TU_INVERT[185]
    '1' & -- TU_INVERT[184]
    '1' & -- TU_INVERT[183]
    '1' & -- TU_INVERT[182]
    '1' & -- TU_INVERT[181]
    '1' & -- TU_INVERT[180]
    '1' & -- TU_INVERT[179]
    '1' & -- TU_INVERT[178]
    '1' & -- TU_INVERT[177]
    '1' & -- TU_INVERT[176]
    '1' & -- TU_INVERT[175]
    '1' & -- TU_INVERT[174]
    '1' & -- TU_INVERT[173]
    '1' & -- TU_INVERT[172]
    '1' & -- TU_INVERT[171]
    '1' & -- TU_INVERT[170]
    '1' & -- TU_INVERT[169]
    '1' & -- TU_INVERT[168]
    '1' & -- TU_INVERT[167]
    '1' & -- TU_INVERT[166]
    '1' & -- TU_INVERT[165]
    '1' & -- TU_INVERT[164]
    '1' & -- TU_INVERT[163]
    '1' & -- TU_INVERT[162]
    '1' & -- TU_INVERT[161]
    '1' & -- TU_INVERT[160]
    '1' & -- TU_INVERT[159]
    '1' & -- TU_INVERT[158]
    '1' & -- TU_INVERT[157]
    '1' & -- TU_INVERT[156]
    '1' & -- TU_INVERT[155]
    '1' & -- TU_INVERT[154]
    '1' & -- TU_INVERT[153]
    '1' & -- TU_INVERT[152]
    '1' & -- TU_INVERT[151]
    '1' & -- TU_INVERT[150]
    '1' & -- TU_INVERT[149]
    '1' & -- TU_INVERT[148]
    '1' & -- TU_INVERT[147]
    '1' & -- TU_INVERT[146]
    '1' & -- TU_INVERT[145]
    '1' & -- TU_INVERT[144]
    '1' & -- TU_INVERT[143]
    '1' & -- TU_INVERT[142]
    '1' & -- TU_INVERT[141]
    '1' & -- TU_INVERT[140]
    '1' & -- TU_INVERT[139]
    '1' & -- TU_INVERT[138]
    '1' & -- TU_INVERT[137]
    '1' & -- TU_INVERT[136]
    '1' & -- TU_INVERT[135]
    '1' & -- TU_INVERT[134]
    '1' & -- TU_INVERT[133]
    '1' & -- TU_INVERT[132]
    '1' & -- TU_INVERT[131]
    '1' & -- TU_INVERT[130]
    '1' & -- TU_INVERT[129]
    '1' & -- TU_INVERT[128]
    '1' & -- TU_INVERT[127]
    '1' & -- TU_INVERT[126]
    '1' & -- TU_INVERT[125]
    '1' & -- TU_INVERT[124]
    '1' & -- TU_INVERT[123]
    '1' & -- TU_INVERT[122]
    '1' & -- TU_INVERT[121]
    '1' & -- TU_INVERT[120]
    '1' & -- TU_INVERT[119]
    '1' & -- TU_INVERT[118]
    '1' & -- TU_INVERT[117]
    '1' & -- TU_INVERT[116]
    '1' & -- TU_INVERT[115]
    '1' & -- TU_INVERT[114]
    '1' & -- TU_INVERT[113]
    '1' & -- TU_INVERT[112]
    '1' & -- TU_INVERT[111]
    '1' & -- TU_INVERT[110]
    '1' & -- TU_INVERT[109]
    '1' & -- TU_INVERT[108]
    '1' & -- TU_INVERT[107]
    '1' & -- TU_INVERT[106]
    '1' & -- TU_INVERT[105]
    '1' & -- TU_INVERT[104]
    '1' & -- TU_INVERT[103]
    '1' & -- TU_INVERT[102]
    '1' & -- TU_INVERT[101]
    '1' & -- TU_INVERT[100]
    '1' & -- TU_INVERT[99]
    '1' & -- TU_INVERT[98]
    '1' & -- TU_INVERT[97]
    '1' & -- TU_INVERT[96]
    '1' & -- TU_INVERT[95]
    '1' & -- TU_INVERT[94]
    '1' & -- TU_INVERT[93]
    '1' & -- TU_INVERT[92]
    '1' & -- TU_INVERT[91]
    '1' & -- TU_INVERT[90]
    '1' & -- TU_INVERT[89]
    '1' & -- TU_INVERT[88]
    '1' & -- TU_INVERT[87]
    '1' & -- TU_INVERT[86]
    '1' & -- TU_INVERT[85]
    '1' & -- TU_INVERT[84]
    '1' & -- TU_INVERT[83]
    '1' & -- TU_INVERT[82]
    '1' & -- TU_INVERT[81]
    '1' & -- TU_INVERT[80]
    '1' & -- TU_INVERT[79]
    '1' & -- TU_INVERT[78]
    '1' & -- TU_INVERT[77]
    '1' & -- TU_INVERT[76]
    '1' & -- TU_INVERT[75]
    '1' & -- TU_INVERT[74]
    '1' & -- TU_INVERT[73]
    '1' & -- TU_INVERT[72]
    '1' & -- TU_INVERT[71]
    '1' & -- TU_INVERT[70]
    '1' & -- TU_INVERT[69]
    '1' & -- TU_INVERT[68]
    '1' & -- TU_INVERT[67]
    '1' & -- TU_INVERT[66]
    '1' & -- TU_INVERT[65]
    '1' & -- TU_INVERT[64]
    '1' & -- TU_INVERT[63]
    '1' & -- TU_INVERT[62]
    '1' & -- TU_INVERT[61]
    '1' & -- TU_INVERT[60]
    '1' & -- TU_INVERT[59]
    '1' & -- TU_INVERT[58]
    '1' & -- TU_INVERT[57]
    '1' & -- TU_INVERT[56]
    '1' & -- TU_INVERT[55]
    '1' & -- TU_INVERT[54]
    '1' & -- TU_INVERT[53]
    '1' & -- TU_INVERT[52]
    '1' & -- TU_INVERT[51]
    '1' & -- TU_INVERT[50]
    '1' & -- TU_INVERT[49]
    '1' & -- TU_INVERT[48]
    '1' & -- TU_INVERT[47]
    '1' & -- TU_INVERT[46]
    '1' & -- TU_INVERT[45]
    '1' & -- TU_INVERT[44]
    '1' & -- TU_INVERT[43]
    '1' & -- TU_INVERT[42]
    '1' & -- TU_INVERT[41]
    '1' & -- TU_INVERT[40]
    '1' & -- TU_INVERT[39]
    '1' & -- TU_INVERT[38]
    '1' & -- TU_INVERT[37]
    '1' & -- TU_INVERT[36]
    '1' & -- TU_INVERT[35]
    '1' & -- TU_INVERT[34]
    '1' & -- TU_INVERT[33]
    '1' & -- TU_INVERT[32]
    '1' & -- TU_INVERT[31]
    '1' & -- TU_INVERT[30]
    '1' & -- TU_INVERT[29]
    '1' & -- TU_INVERT[28]
    '1' & -- TU_INVERT[27]
    '1' & -- TU_INVERT[26]
    '1' & -- TU_INVERT[25]
    '1' & -- TU_INVERT[24]
    '1' & -- TU_INVERT[23]
    '1' & -- TU_INVERT[22]
    '1' & -- TU_INVERT[21]
    '1' & -- TU_INVERT[20]
    '1' & -- TU_INVERT[19]
    '1' & -- TU_INVERT[18]
    '1' & -- TU_INVERT[17]
    '1' & -- TU_INVERT[16]
    '1' & -- TU_INVERT[15]
    '1' & -- TU_INVERT[14]
    '1' & -- TU_INVERT[13]
    '1' & -- TU_INVERT[12]
    '1' & -- TU_INVERT[11]
    '1' & -- TU_INVERT[10]
    '1' & -- TU_INVERT[9]
    '1' & -- TU_INVERT[8]
    '1' & -- TU_INVERT[7]
    '1' & -- TU_INVERT[6]
    '1' & -- TU_INVERT[5]
    '1' & -- TU_INVERT[4]
    '1' & -- TU_INVERT[3]
    '1' & -- TU_INVERT[2]
    '1' & -- TU_INVERT[1]
    '1' ; -- TU_INVERT[0]

end package;
