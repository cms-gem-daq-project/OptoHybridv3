----------------------------------------------------------------------------------
-- CMS Muon Endcap
-- GEM Collaboration
-- Optohybrid v3 Firmware -- Clocking
-- 2017/07/21 -- Initial port to version 3 electronics
-- 2017/07/22 -- Additional MMCM added to monitor and dejitter the eport clock
-- 2017/08/09 -- 200MHz iodelay refclk added to primary MMCM
-- 2019/05/02 -- Added BUFGCE outputs to disable clocks during MGT init
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

library work;
use work.types_pkg.all;
use work.param_pkg.all;
use work.ipbus_pkg.all;
use work.registers.all;

entity clocking is
generic(
    g_ERROR_COUNT_MAX : integer := 5;
    g_DONT_USE_CLOCK_GATING : std_logic := '0'
);
port(

    clock_p : in std_logic;
    clock_n : in std_logic;

    clk40_o      : out std_logic; -- 40 MHz phase shiftable frame clock from GBT
    clk80_o      : out std_logic; -- 80 MHz phase shiftable frame clock from GBT
    clk160_0_o   : out std_logic; -- 160 MHz phase shiftable frame clock from GBT
    clk160_90_o  : out std_logic; -- 160 MHz phase shiftable frame clock from GBT
    clk200_o     : out std_logic;

    -- mmcm locked status monitors
    mmcm_locked_o   : out std_logic;

    -- ipbus

    ipb_mosi_i : in  ipb_wbus;
    ipb_miso_o : out ipb_rbus;

    ipb_reset_i : in std_logic;

    cnt_snap : in std_logic

);
end clocking;


architecture Behavioral of clocking is

    signal clk40      : std_logic; -- 40 MHz phase shiftable frame clock from GBT
    signal clk80      : std_logic; -- 80 MHz phase shiftable frame clock from GBT
    signal clk160_0   : std_logic; -- 160 MHz phase shiftable frame clock from GBT
    signal clk160_90  : std_logic; -- 160 MHz phase shiftable frame clock from GBT
    signal clk200     : std_logic;

    signal mmcm_locked : std_logic;

    signal clock   : std_logic;
    signal clock_i : std_logic;

    ------ Register signals begin (this section is generated by <optohybrid_top>/tools/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_write_arr       : t_std32_array(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_addresses       : t_std32_array(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_defaults        : t_std32_array(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => '0');
    signal regs_write_pulse_arr : std_logic_vector(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => '0');
    signal regs_read_ready_arr  : std_logic_vector(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_CLOCKING_NUM_REGS - 1 downto 0) := (others => '0');
    -- Connect counter signal declarations
    signal mmcm_unlocked : std_logic_vector (7 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------

begin

      -- Input buffering
      --------------------------------------
    clkin1_buf : IBUFGDS
    port map (
        O  => clock_i,
        I  => clock_p,
        IB => clock_n
    );

    logic_clocking : entity work.logic_clocking
    port map(

        clk_in1     => clock_i,

        clk40_o     => clk40,
        clk80_o     => clk80,
        clk160_o    => clk160_0,
        clk160_90_o => clk160_90,
        clk200_o    => clk200,

        locked_o    => mmcm_locked
    );

    clk40_o      <=     clk40;
    clk80_o      <=     clk80;
    clk160_0_o   <=     clk160_0;
    clk160_90_o  <=     clk160_90;
    clk200_o     <=     clk200;

    mmcm_locked_o <= mmcm_locked;

    --===============================================================================================
    -- (this section is generated by <optohybrid_top>/tools/generate_registers.py -- do not edit)
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_CLOCKING_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_CLOCKING_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_CLOCKING_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => clock,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => clock,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_CLOCKING_ADDRESS_MSB downto REG_CLOCKING_ADDRESS_LSB) <= "00";

    -- Connect read signals
    regs_read_arr(0)(REG_CLOCKING_MMCM_LOCKED_BIT) <= mmcm_locked;
    regs_read_arr(0)(REG_CLOCKING_MMCM_UNLOCKED_CNT_MSB downto REG_CLOCKING_MMCM_UNLOCKED_CNT_LSB) <= mmcm_unlocked;

    -- Connect write signals

    -- Connect write pulse signals

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect counter instances

    COUNTER_CLOCKING_MMCM_UNLOCKED_CNT : entity work.counter_snap
    generic map (
        g_COUNTER_WIDTH  => 8
    )
    port map (
        ref_clk_i => clock,
        reset_i   => ipb_reset_i,
        en_i      => not mmcm_locked,
        snap_i    => '1',
        count_o   => mmcm_unlocked
    );


    -- Connect rate instances

    -- Connect read ready signals

    -- Defaults

    -- Define writable regs

    --==== Registers end ============================================================================

end Behavioral;
